//import "DPI-C" function string getenv(input string env_name);

module top_tb;

    timeunit 1ps;
    timeprecision 1ps;

    //int clock_half_period_ps = getenv("ECE411_CLOCK_PERIOD_PS").atoi() / 2;
    int clock_half_period_ps = 10 / 2;

    bit clk;
    always #(clock_half_period_ps) clk = ~clk;

    bit rst;

    int timeout = 10000000; // in cycles, change according to your needs


    mem_itf_banked bmem_itf(.*);

   `ifdef RND_TEST
    random_tb random_tb(.itf(bmem_itf)); // For randomized testing
    rob_mon  rob_tom ( .* , .rob2mon_itf( dut.u_ooo.rob2mon_itf ) ) ;
    `else
    banked_memory banked_memory(.itf(bmem_itf));
    `endif

    mon_itf #(.CHANNELS(8)) mon_itf(.*);
    monitor #(.CHANNELS(8)) monitor(.itf(mon_itf));

    cpu dut(
        .clk            (clk),
        .rst            (rst),

        .bmem_addr  (bmem_itf.addr  ),
        .bmem_read  (bmem_itf.read  ),
        .bmem_write (bmem_itf.write ),
        .bmem_wdata (bmem_itf.wdata ),
        .bmem_ready (bmem_itf.ready ),
        .bmem_raddr (bmem_itf.raddr ),
        .bmem_rdata (bmem_itf.rdata ),
        .bmem_rvalid(bmem_itf.rvalid)
    );

    `include "rvfi_reference.svh"

    initial begin
        $fsdbDumpfile("dump.fsdb");
        $fsdbDumpvars(0, "+all");
        rst = 1'b1;
        repeat (2) @(posedge clk);
        rst <= 1'b0;

    end

    always @(posedge clk) begin
        for (int unsigned i=0; i < 8; ++i) begin
            if (mon_itf.halt[i]) begin
                $finish;
            end
        end
        if (timeout == 0) begin
            $error("TB Error: Timed out");
            $finish;
        end
        if (mon_itf.error != 0) begin
            repeat (15) @(posedge clk);
            $finish;
        end
        if (bmem_itf.error != 0) begin
            repeat (5) @(posedge clk);
            $finish;
        end
        timeout <= timeout - 1;
    end

endmodule
